-- Testbench for 74154 TTL demultiplexer
library IEEE;
use IEEE.std_logic_1164.all;
 
entity testbench is
-- empty
end testbench; 

architecture tb of testbench is

-- DUT component

component TTL74154 is
port(
  pin1_ny0  : out std_logic;
  pin2_ny1  : out std_logic;
  pin3_ny2  : out std_logic;
  pin4_ny3  : out std_logic;
  pin5_ny4  : out std_logic;
  pin6_ny5  : out std_logic;
  pin7_ny6  : out std_logic;
  pin8_ny7  : out std_logic;
  pin9_ny8  : out std_logic;
  pin10_ny9  : out std_logic;
  pin11_ny10  : out std_logic;  
  pin13_ny11  : out std_logic;
  pin14_ny12  : out std_logic;
  pin15_ny13  : out std_logic;
  pin16_ny14: out std_logic;
  pin17_ny15: out std_logic;  
  pin18_ne1: in std_logic;
  pin19_ne2: in std_logic;
  pin20_a3: in std_logic;
  pin21_a2: in std_logic;
  pin22_a1 : in std_logic;
  pin23_a0 : in std_logic);
end component;

signal ny0,ny1,ny2,ny3,ny4,ny5,ny6,ny7,ny8,ny9,ny10,ny11,ny12,ny13,ny14,ny15,ne1,ne2,a3,a2,a1,a0: std_logic;
begin

  -- Connect DUT
  DUT: TTL74154 port map(ny0,ny1,ny2,ny3,ny4,ny5,ny6,ny7,ny8,ny9,ny10,ny11,ny12,ny13,ny14,ny15,ne1,ne2,a3,a2,a1,a0);
  process
  begin
    ne1 <= '1';
    ne2 <= '1';
    a3 <= 'X';
    a2 <= 'X';
    a1 <= 'X';
    a0 <= 'X';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;

    ne1 <= '0';
    ne2 <= '1';
    a3 <= 'X';
    a2 <= 'X';
    a1 <= 'X';
    a0 <= 'X';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '1';
    ne2 <= '0';
    a3 <= 'X';
    a2 <= 'X';
    a1 <= 'X';
    a0 <= 'X';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;

    ne1 <= '0';
    ne2 <= '0';
    a3 <= '0';
    a2 <= '0';
    a1 <= '0';
    a0 <= '0';
    wait for 100 ns;
    assert (ny0 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '0';
    a2 <= '0';
    a1 <= '0';
    a0 <= '1';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '0';
    a2 <= '0';
    a1 <= '1';
    a0 <= '0';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '0';
    a2 <= '0';
    a1 <= '1';
    a0 <= '1';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '0';
    a2 <= '1';
    a1 <= '0';
    a0 <= '0';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '0';
    a2 <= '1';
    a1 <= '0';
    a0 <= '1';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '0';
    a2 <= '1';
    a1 <= '1';
    a0 <= '0';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '0';
    a2 <= '1';
    a1 <= '1';
    a0 <= '1';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '1';
    a2 <= '0';
    a1 <= '0';
    a0 <= '0';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '1';
    a2 <= '0';
    a1 <= '0';
    a0 <= '1';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;

    ne1 <= '0';
    ne2 <= '0';
    a3 <= '1';
    a2 <= '0';
    a1 <= '1';
    a0 <= '0';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
 
 
     ne1 <= '0';
    ne2 <= '0';
    a3 <= '1';
    a2 <= '0';
    a1 <= '1';
    a0 <= '1';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '1';
    a2 <= '1';
    a1 <= '0';
    a0 <= '0';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny1 not set" severity error;
    assert (ny2 = '1') report "Fail ny2 not set" severity error;
    assert (ny3 = '1') report "Fail ny3 not set" severity error;
    assert (ny4 = '1') report "Fail ny4 not set" severity error;
    assert (ny5 = '1') report "Fail ny5 not set" severity error;
    assert (ny6 = '1') report "Fail ny6 not set" severity error;
    assert (ny7 = '1') report "Fail ny7 not set" severity error;
    assert (ny8 = '1') report "Fail ny8 not set" severity error;
    assert (ny9 = '1') report "Fail ny9 not set" severity error;
    assert (ny10 = '1') report "Fail ny10 not set" severity error;
    assert (ny11 = '1') report "Fail ny11 not set" severity error;
    assert (ny12 = '0') report "Fail ny12 not cleared" severity error;
    assert (ny13 = '1') report "Fail ny13 not set" severity error;
    assert (ny14 = '1') report "Fail ny14 not set" severity error;
    assert (ny15 = '1') report "Fail ny15 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '1';
    a2 <= '1';
    a1 <= '0';
    a0 <= '1';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '1';
    a2 <= '1';
    a1 <= '1';
    a0 <= '0';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '0') report "Fail ny0 not cleared" severity error;
    assert (ny15 = '1') report "Fail ny0 not set" severity error;
    
    ne1 <= '0';
    ne2 <= '0';
    a3 <= '1';
    a2 <= '1';
    a1 <= '1';
    a0 <= '1';
    wait for 100 ns;
    assert (ny0 = '1') report "Fail ny0 not set" severity error;
    assert (ny1 = '1') report "Fail ny0 not set" severity error;
    assert (ny2 = '1') report "Fail ny0 not set" severity error;
    assert (ny3 = '1') report "Fail ny0 not set" severity error;
    assert (ny4 = '1') report "Fail ny0 not set" severity error;
    assert (ny5 = '1') report "Fail ny0 not set" severity error;
    assert (ny6 = '1') report "Fail ny0 not set" severity error;
    assert (ny7 = '1') report "Fail ny0 not set" severity error;
    assert (ny8 = '1') report "Fail ny0 not set" severity error;
    assert (ny9 = '1') report "Fail ny0 not set" severity error;
    assert (ny10 = '1') report "Fail ny0 not set" severity error;
    assert (ny11 = '1') report "Fail ny0 not set" severity error;
    assert (ny12 = '1') report "Fail ny0 not set" severity error;
    assert (ny13 = '1') report "Fail ny0 not set" severity error;
    assert (ny14 = '1') report "Fail ny0 not set" severity error;
    assert (ny15 = '0') report "Fail ny0 not cleared" severity error;    
    
	assert false report "Test done." severity note;
    wait;
  end process;
end tb;

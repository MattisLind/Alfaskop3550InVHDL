-- Testbench for 74193 TTL counter
library IEEE;
use IEEE.std_logic_1164.all;
 
entity testbench is
-- empty
end testbench; 

architecture tb of testbench is

-- DUT component

component TTL74193 is
port(
  pin1_b  : in std_logic;
  pin2_qB   : out std_logic;
  pin3_qA   : out std_logic;
  pin4_down: in std_logic;
  pin5_up  : in std_logic;
  pin6_qC   : out std_logic;
  pin7_qD   : out std_logic;
  pin9_d  : in std_logic;
  pin10_c : in std_logic;
  pin11_nLoad: in std_logic;  
  pin12_nCO : out std_logic;
  pin13_nBO : out std_logic;
  pin14_clr: in std_logic;
  pin15_a : in std_logic);
end component;

signal b,qB,qA,down,up,qC,qD,d,c,nLoad,nCO,nBO,clr,a: std_logic;
begin

  -- Connect DUT
  DUT: TTL74193 port map(b,qB,qA,down,up,qC,qD,d,c,nLoad,nCO,nBO,clr,a);
  process
  begin
    a <= '0';
    b <= '0';
    c <='0';
    d <= '0';
    up <= '1';
    down <='1';
    nLoad <= '1';
    clr <= '0';
    wait for 100 ns;
    clr <= '1';
    wait for 100 ns;
    clr <= '0';
	assert (qA = '0') report "Fail qA not cleared" severity error;
    assert (qB = '0') report "Fail qB not cleared" severity error;
    assert (qC = '0') report "Fail qC not cleared" severity error;
    assert (qD = '0') report "Fail qD not cleared" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    a  <= '1';
    b  <= '0';
    c  <= '0';
    d  <= '1';
    nLoad <= '0';
    wait for 100 ns;
    nLoad <= '1';
    assert (qA = '1') report "Fail qA not set after load" severity error;
    assert (qB = '0') report "Fail qB not cleared after load" severity error;
    assert (qC = '0') report "Fail qC not cleared after load" severity error;
    assert (qD = '1') report "Fail qD not set after load" severity error;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    up <= '0';
    wait for 100 ns;
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '0') report "Fail qA not cleared after count up" severity error;
    assert (qB = '1') report "Fail qB not set after count up" severity error;
    assert (qC = '0') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;    
    up <= '0';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '1') report "Fail qA not set after count up" severity error;
    assert (qB = '1') report "Fail qB not set after count up" severity error;
    assert (qC = '0') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;
    up <= '0';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nCO not set after count up" severity error;
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '0') report "Fail qA not set after count up" severity error;
    assert (qB = '0') report "Fail qB not set after count up" severity error;
    assert (qC = '1') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;
    up <= '0';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nCO not set after count up" severity error;
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '1') report "Fail qA not set after count up" severity error;
    assert (qB = '0') report "Fail qB not set after count up" severity error;
    assert (qC = '1') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;
    up <= '0';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '0') report "Fail qA not set after count up" severity error;
    assert (qB = '1') report "Fail qB not set after count up" severity error;
    assert (qC = '1') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;
    up <= '0';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '1') report "Fail qA not set after count up" severity error;
    assert (qB = '1') report "Fail qB not set after count up" severity error;
    assert (qC = '1') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;    
    up <= '0';
    wait for 100 ns;
    assert (nCO = '0') report "Fail nCO not cleared after count up to carry" severity error; 
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '0') report "Fail qA not set after count up" severity error;
    assert (qB = '0') report "Fail qB not set after count up" severity error;
    assert (qC = '0') report "Fail qC not cleared after count up" severity error;
    assert (qD = '0') report "Fail qD not set after count up" severity error;    
    up <= '0';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not cleared after count up to carry" severity error; 
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '1') report "Fail qA not set after count up" severity error;
    assert (qB = '0') report "Fail qB not set after count up" severity error;
    assert (qC = '0') report "Fail qC not cleared after count up" severity error;
    assert (qD = '0') report "Fail qD not set after count up" severity error;    
    up <= '0';
    wait for 100 ns;
    assert (nBO = '1') report "Fail nCO not set after count up" severity error;
    assert (nCO = '1') report "Fail nBO not cleared after count up to carry" severity error;  
    up <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '0') report "Fail qA not set after count up" severity error;
    assert (qB = '1') report "Fail qB not set after count up" severity error;
    assert (qC = '0') report "Fail qC not cleared after count up" severity error;
    assert (qD = '0') report "Fail qD not set after count up" severity error;    
    down <= '0';
    wait for 100 ns;
    assert (nBO = '1') report "Fail nCO not set after count up" severity error;
    assert (nCO = '1') report "Fail nCO not cleared after count up to carry" severity error; 
    down <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '1') report "Fail qA not set after count up" severity error;
    assert (qB = '0') report "Fail qB not set after count up" severity error;
    assert (qC = '0') report "Fail qC not cleared after count up" severity error;
    assert (qD = '0') report "Fail qD not set after count up" severity error;
    down <= '0';
    wait for 100 ns;
    assert (nBO = '1') report "Fail nCO not set after count up" severity error;
    assert (nCO = '1') report "Fail nCO not cleared after count up to carry" severity error; 
    down <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '0') report "Fail qA not set after count up" severity error;
    assert (qB = '0') report "Fail qB not set after count up" severity error;
    assert (qC = '0') report "Fail qC not cleared after count up" severity error;
    assert (qD = '0') report "Fail qD not set after count up" severity error;
    down <= '0';
    wait for 100 ns;
    assert (nBO = '0') report "Fail nCO not set after count up" severity error;
    assert (nCO = '1') report "Fail nCO not cleared after count up to carry" severity error; 
    down <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '1') report "Fail qA not set after count up" severity error;
    assert (qB = '1') report "Fail qB not set after count up" severity error;
    assert (qC = '1') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;
    down <= '0';
    wait for 100 ns;
    assert (nBO = '1') report "Fail nCO not set after count up" severity error;
    assert (nCO = '1') report "Fail nCO not cleared after count up to carry" severity error; 
    down <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '0') report "Fail qA not set after count up" severity error;
    assert (qB = '1') report "Fail qB not set after count up" severity error;
    assert (qC = '1') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;
    down <= '0';
    wait for 100 ns;
    assert (nBO = '1') report "Fail nCO not set after count up" severity error;
    assert (nCO = '1') report "Fail nCO not cleared after count up to carry" severity error; 
    down <= '1';
    wait for 100 ns;
    assert (nCO = '1') report "Fail nCO not set after count up" severity error;
    assert (nBO = '1') report "Fail nBO not set after count up" severity error;
    assert (qA = '1') report "Fail qA not set after count up" severity error;
    assert (qB = '0') report "Fail qB not set after count up" severity error;
    assert (qC = '1') report "Fail qC not cleared after count up" severity error;
    assert (qD = '1') report "Fail qD not set after count up" severity error;    
	assert false report "Test done." severity note;
    wait;
  end process;
end tb;

-- Testbench for 74198 TTL shift register
library IEEE;
use IEEE.std_logic_1164.all;
 
entity testbench is
-- empty
end testbench; 

architecture tb of testbench is

-- DUT component

component TTL74198 is
port(
  pin1_s0: in std_logic;
  pin2_srsi  : in std_logic;
  pin3_a : in std_logic;
  pin4_qA   : out std_logic;
  pin5_b  : in std_logic;
  pin6_qB   : out std_logic;
  pin7_c : in std_logic;
  pin8_qC   : out std_logic;
  pin9_d  : in std_logic;
  pin10_qD   : out std_logic;
  pin11_clk: in std_logic;
  pin13_clear : in std_logic;
  pin14_qE   : out std_logic;
  pin15_e : in std_logic;
  pin16_qF   : out std_logic;
  pin17_f  : in std_logic;
  pin18_qG   : out std_logic;
  pin19_g : in std_logic;
  pin20_qH   : out std_logic;
  pin21_h  : in std_logic;
  pin22_slsi : in std_logic;
  pin23_s1: in std_logic);
end component;

signal s0,srsi,a,qA,b,qB,c,qC,d,qD,clk,clear,qE,e,qF,f,qG,g,qH,h,slsi,s1: std_logic;
begin

  -- Connect DUT
  DUT: TTL74198 port map(s0,srsi,a,qA,b,qB,c,qC,d,qD,clk,clear,qE,e,qF,f,qG,g,qH,h,slsi,s1);
  process
  begin
    clk <= '0';
    srsi <= '0';
    s0 <='0';
    s1 <= '0';
    a <= '0';
    b <= '0';
    c <= '0';
    d <= '0';
    e <= '0';
    f <= '0';
    g <= '0';
    h <= '0';
    slsi <= '0';
    clear <= '0';
    wait for 100 ns;
	assert (qA = '0') report "Fail qA not cleared" severity error;
    assert (qB = '0') report "Fail qB not cleared" severity error;
    assert (qC = '0') report "Fail qC not cleared" severity error;
    assert (qD = '0') report "Fail qD not cleared" severity error;
	assert (qE = '0') report "Fail qE not cleared" severity error;
    assert (qF = '0') report "Fail qF not cleared" severity error;
    assert (qG = '0') report "Fail qG not cleared" severity error;
    assert (qH = '0') report "Fail qH not cleared" severity error;
    clear <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not cleared" severity error;
    assert (qB = '0') report "Fail qB not cleared" severity error;
    assert (qC = '0') report "Fail qC not cleared" severity error;
    assert (qD = '0') report "Fail qD not cleared" severity error;
	assert (qE = '0') report "Fail qE not cleared" severity error;
    assert (qF = '0') report "Fail qF not cleared" severity error;
    assert (qG = '0') report "Fail qG not cleared" severity error;
    assert (qH = '0') report "Fail qH not cleared" severity error;
    a  <= '1';
    b  <= '0';
    c  <= '1';
    d  <= '0';
    e  <= '1';
    f  <= '0';
    g  <= '1';
    h  <= '1';
    s0 <= '1';
    s1 <= '1';
	wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '1') report "Fail qA not loaded" severity error;
    assert (qB = '0') report "Fail qB not loaded" severity error;
    assert (qC = '1') report "Fail qC not loaded" severity error;
    assert (qD = '0') report "Fail qD not loaded" severity error;
	assert (qE = '1') report "Fail qE not loaded" severity error;
    assert (qF = '0') report "Fail qF not loaded" severity error;
    assert (qG = '1') report "Fail qG not loaded" severity error;
    assert (qH = '1') report "Fail qH not loaded" severity error;
    clk <= '0';
    wait for 100 ns;
    assert (qA = '1') report "Fail qA not loaded" severity error;
    assert (qB = '0') report "Fail qB not loaded" severity error;
    assert (qC = '1') report "Fail qC not loaded" severity error;
    assert (qD = '0') report "Fail qD not loaded" severity error;
	assert (qE = '1') report "Fail qE not loaded" severity error;
    assert (qF = '0') report "Fail qF not loaded" severity error;
    assert (qG = '1') report "Fail qG not loaded" severity error;
    assert (qH = '1') report "Fail qH not loaded" severity error;
    s0 <= '1';
    s1 <= '0';
    srsi <= '0';
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '1') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error;
	clk <= '0';
    wait for 100 ns;
    srsi <= '1';
    clk <= '1';
    wait for 100 ns;
    assert (qA = '1') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '1') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '1') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '1') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error;
    clk <= '0';
    wait for 100 ns;
    srsi <= '0';
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '1') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error;
    clk <= '0';
    wait for 100 ns;
    srsi <= '0';
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '1') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '1') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '1') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error;
    clk <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error;
    clk <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '1') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '1') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error;   
    clk <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error;    
    clk <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '1') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error;   
    clk <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error;   
    clk <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error; 
    wait for 100 ns;
    s0 <= '0';
    s1 <= '1';
    wait for 100 ns;
    clk <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error; 
    clk <= '0';
    slsi <= '1';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    clk <= '0';
    slsi <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '1') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error; 
    clk <= '0';
    slsi <= '1';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    clk <= '0';
    slsi <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '1') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '1') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error; 
    clk <= '0';
    slsi <= '1';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    clk <= '0';
    slsi <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '1') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '1') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '1') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error; 
    clk <= '0';
    slsi <= '1';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '1') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    wait for 100 ns;
	s1 <= '0';	
    clk <= '0';
    slsi <= '1';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '1') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    wait for 100 ns;
	s1 <= '0';	
    clk <= '0';
    slsi <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '1') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    wait for 100 ns;
	s1 <= '0';	
    clk <= '0';
    slsi <= '1';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '1') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    wait for 100 ns;
	s1 <= '0';	
    clk <= '0';
    slsi <= '0';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '1') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    wait for 100 ns;
    clk <= '0';
    slsi <= '1';
    wait for 100 ns;
    clk <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '1') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '1') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '1') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '1') report "Fail qH not shifted in" severity error; 
    wait for 100 ns;
	clear <= '0';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error; 
    wait for 100 ns;
	clear <= '1';
    wait for 100 ns;
    assert (qA = '0') report "Fail qA not shifted in" severity error;
    assert (qB = '0') report "Fail qB not shifted in" severity error;
    assert (qC = '0') report "Fail qC not shifted in" severity error;
    assert (qD = '0') report "Fail qD not shifted in" severity error;    
	assert (qE = '0') report "Fail qE not shifted in" severity error;
    assert (qF = '0') report "Fail qF not shifted in" severity error;
    assert (qG = '0') report "Fail qG not shifted in" severity error;
    assert (qH = '0') report "Fail qH not shifted in" severity error; 
    
	assert false report "Test done." severity note;
    wait;
  end process;
end tb;
